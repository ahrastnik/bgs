library IEEE;
use IEEE.numeric_std.all;
use IEEE.std_logic_1164.all;

entity GPU is
	port(
		clk: in std_logic
	);
end GPU;

architecture Malibu of GPU is
	
begin
	
end Malibu;